the 149 of 111 to 91 and 87 I 76 my 55 a 50 in 41 was 35 that 33 had 33 but 24 his 22 have 21 which 21 me 19 not 19 her 19 were 17 with 17 as 16 at 13 for 12 been 12 He 11 from 11 he 11 M. 10 is 10 it 10 be 10 by 10 natural 9 she 9 you 9 on 9 your 9 when 9 She 8 one 8 those 8 The 7 these 7 upon 7 science 7 own 7 an 7 My 6 this 6 they 6 day 6 modern 6 new 6 said 6 we 6 whom 6 life 6 myself 6 into 6 made 6 other 6 father 5 very 5 little 5 would 5 must 5 can 5 so 5 Elizabeth 5 first 5 most 5 should 5 are 5 will 5 concerning 5 whose 4 persuade 4 even 4 professor 4 studies 4 names 4 rather 4 its 4 then 4 now 4 given 4 could 4 such 4 spent 4 Krempe 4 reflections 4 during 4 fellow 4 It 4 greatest 4 They 4 some 4 or 4 lecture 4 books 4 no 4 time 4 all 3 more, 3 did 3 what 3 principal 3 ever 3 never 3 desired 3 same 3 more 3 grief 3 account 3 said, 3 different 3 man 3 departure 3 over 3 His 3 our 3 attended 3 length 3 their 3 Such 3 than 3 youth 3 Waldman, 3 any 3 hitherto 3 philosophy 3 took 3 future 3 science. 3 only 3 men 3 away 3 various 3 many 3 appeared 3 ourselves 3 voice 3 itself 3 In 3 if 3 thought 3 without 3 mother 3 has 3 ought 3 On 3 world 3 steps 3 become 3 dear 3 felt 3 although 3 after 3 long 3 Ingolstadt, 3 philosophy. 3 remarkably 2 And 2 returned 2 went 2 list 2 her. 2 me, 2 me. 2 me; 2 deeply 2 expressed 2 degree 2 eye 2 few 2 ambition 2 So 2 age, 2 us. 2 soul 2 believed 2 heard 2 heard. 2 performed 2 contempt 2 how 2 intended 2 may 2 chiefly 2 every 2 nearly 2 replied 2 indeed 2 soon 2 years 2 course 2 before 2 them 2 evening 2 hands 2 masters 2 university 2 each 2 entirely 2 house 2 hard 2 out 2 misfortune 2 time, 2 attentions 2 This 2 bestow 2 Waldman 2 days 2 place 2 improvements 2 Elizabeth, 2 ancient 2 eyes 2 authors 2 branches 2 morning's 2 illness 2 remained 2 mind 2 say 2 rent 2 saw 2 paid 2 connected 2 alone. 2 hopes 2 chord 2 We 2 knowledge 2 state 2 repose, 2 familiar 2 words 2 him 2 enough 2 nature 2 regret 2 last 2 gave 2 quit 2 But 2 duties 2 partly 2 make 2 several 2 week 2 hand 2 uses 2 thoughts 2 chemistry 2 being 2 human 2 beloved 2 useless 2 resolved 2 explained 2 early 2 acquainted 2 delivered 2 Clerval 2 there 2 us 2 convey 2 describe 2 am 2 knowledge. 2 again 2 branch 2 evil, 2 desert 2 As 2 far 2  1 results 1 son. 1 reflections. 1 mild 1 burdened 1 benevolence; 1 go 1 directed, 1 fatiguing. 1 reluctant 1 devoted 1 acquired 1 apartment 1 fancies 1 steadily 1 presents 1 present 1 under 1 smile 1 sorry 1 fatal 1 sway 1 advantage 1 void 1 (inexperience 1 strangers. 1 "every 1 soul, 1 worst 1 presumption 1 Henry 1 classifications 1 continued 1 recollected 1 treating 1 discovered 1 joined 1 leave 1 solid 1 retrod 1 steeple 1 circulates, 1 concluded 1 lecturing 1 among 1 playmate 1 children," 1 air 1 expressive 1 saved, 1 prepossess 1 plays 1 town. 1 calmly, 1 Clerval; 1 seen, 1 musty 1 ended 1 above 1 entreaties, 1 During 1 filled 1 deemed 1 led 1 exchange 1 doubt 1 hairs 1 equals 1 explore 1 made; 1 let 1 conceited 1 along 1 extreme 1 obtained 1 great 1 animated 1 statement, 1 professors. 1 light. 1 banished. 1 elixir 1 discoveries 1 women 1 descended 1 permit 1 residents 1 unknown 1 consoled. 1 felt, 1 consolation 1 thought, 1 sweetest 1 merely 1 world." 1 When 1 private 1 feelings 1 ascend 1 relations, 1 deceived; 1 science," 1 glance 1 "my 1 public, 1 use 1 spoke 1 remains 1 Agrippa 1 visit 1 two 1 next 1 going 1 call 1 therefore 1 memory 1 taken 1 misery. 1 God! 1 gained 1 door 1 befitting 1 These 1 idleness, 1 company 1 Krempe, 1 occurred 1 refrain 1 sorrow, 1 commenced 1 ardently 1 awoke, 1 former 1 debarred 1 foundations 1 "to 1 task, 1 and, 1 Now 1 word 1 lapse 1 us, 1 gruff 1 remain 1 irreparable 1 learn 1 akin 1 shadows." 1 nothing. 1 degrees, 1 requested, 1 history 1 control 1 indulgence 1 "old 1 give 1 neglected 1 high 1 want 1 sought 1 cursory 1 native 1 information 1 labours. 1 grand; 1 renew 1 dismissed 1 fortunate 1 write 1 kindness. 1 extinguished 1 alighted 1 mysteries 1 "My 1 A 1 fever 1 rude 1 advice 1 act 1 genius, 1 customs 1 purpose. 1 produce 1 strove 1 blood 1 curiosity 1 ties 1 journey; 1 short 1 third 1 discoverers. 1 endeavoured 1 exhibited 1 inform 1 cannot 1 enter 1 procure. 1 procure, 1 learning, 1 began 1 modesty 1 would, 1 devote 1 exclaimed 1 countenances. 1 professors 1 ashamed) 1 dearest 1 including 1 looks 1 affectation, 1 penetrate 1 mentioned 1 existence 1 still 1 solitary 1 thence 1 bringing 1 labours 1 stimulated 1 immortality 1 systems 1 dead, 1 covered 1 arrange 1 easier 1 I, 1 it. 1 return 1 little, 1 indefatigable 1 sounded, 1 professor. 1 prejudices 1 professor, 1 little; 1 repulsive 1 nor 1 possess 1 came. 1 brightness 1 all. 1 all, 1 whither 1 creation. 1 bless 1 tear 1 sleep 1 all? 1 accompanied 1 happy," 1 met 1 pursuits 1 disciple; 1 elementary 1 therefore, 1 taught 1 forgot 1 dawn 1 indulged 1 "really 1 alchemists. 1 surrounded 1 futile, 1 keys 1 boundless 1 inquirer 1 Frankenstein 1 fortitude 1 pulpit, 1 appertaining 1 turning 1 mourning 1 attending 1 alchemists 1 enlightened 1 beginning 1 ability, 1 pursuits. 1 perhaps, 1 fever; 1 due 1 After 1 domestic, 1 conducted 1 black. 1 think 1 perform; 1 mathematics." 1 indebted 1 already 1 peculiar 1 stared. 1 anxiety. 1 There 1 brothers, 1 philosophical 1 "Farewell!" 1 another 1 comforter 1 thick 1 thousand 1 reprobated; 1 cheerfully 1 introduction 1 love, 1 caught 1 station 1 power; 1 too 1 white 1 recent 1 really 1 colleague. 1 attendants 1 mentioning 1 accompany 1 exploded 1 changed. 1 part 1 forget: 1 wasted 1 herself 1 sickened; 1 spoiler 1 kind 1 hushed, 1 night. 1 folly 1 views, 1 bitterness 1 omitted. 1 upon. 1 chemists; 1 miracles. 1 distinguished 1 acquisition 1 prospect 1 recesses 1 sentences 1 need 1 Albertus 1 sat 1 paths 1 squat 1 narrow-minded 1 thunders 1 general 1 studying 1 often, 1 uncouth 1 aside 1 distemper 1 localities 1 breathe. 1 take 1 late. 1 chaise 1 With 1 lectures 1 begin 1 added 1 amiable 1 shall 1 countenance. 1 machines, 1 Good 1 pleasure 1 Partly 1 measured 1 why 1 sickbed; 1 spirits 1 forever 1 consequences 1 feminine 1 considered 1 medical 1 panegyric 1 order 1 looked 1 accounted 1 terms, 1 uncle 1 If 1 promising 1 saying, 1 lived, 1 terms. 1 show 1 favour 1 fervour 1 companions, 1 "These 1 find 1 feel? 1 arrived. 1 completion 1 with, 1 founded. 1 advanced 1 abode. 1 ruin 1 cousins. 1 sacrilege 1 erect 1 touched 1 pretty 1 consent 1 attained 1 chemistry, 1 entreaties 1 hope 1 exchanged 1 heaven, 1 closed 1 listened 1 loved 1 kindling 1 leave. 1 enemy; 1 expectation 1 leisure 1 yielded 1 courage 1 weeks. 1 warmth, 1 crucible, 1 commerce. 1 way, 1 following 1 resolve 1 scene 1 Angel 1 whilst 1 seemed 1 command 1 affability 1 heavens; 1 morning 1 "Every 1 microscope 1 wish 1 fixed 1 where 1 wrote 1 beings. 1 seventeen 1 questions 1 triumphed 1 melancholy 1 mechanism 1 symptoms, 1 grey 1 see 1 decided 1 hear 1 fail 1 miserable 1 best 1 powers, 1 annihilation 1 repugnance 1 matters, 1 mien 1 aspirations 1 alarming 1 firmest 1 protector. 1 strain, 1 continually 1 father's 1 determined 1 years. 1 progress 1 man, 1 date, 1 faces," 1 terms 1 days; 1 commence 1 confusion 1 sorrow 1 attention 1 deliver 1 sacrilege, 1 however 1 countenance 1 Thus 1 unfold 1 invisible 1 dawn, 1 connection? 1 proceeded, 1 influence, 1 repent. 1 secrets 1 trader 1 escape 1 powers; 1 against 1 union. 1 forgotten 1 Cornelius 1 Yet 1 journey 1 supply 1 sweet 1 aspect 1 manners 1 achieve; 1 asserted 1 complied 1 arise, 1 petty 1 recur 1 come 1 teacher, 1 three 1 were, 1 Chance 1 experiments, 1 philosophers, 1 interest 1 entered 1 meeting 1 instructing 1 threw 1 firm 1 success. 1 turned 1 sufficient 1 sunshine 1 imprudence 1 recalled 1 child 1 instant 1 realities 1 sound 1 yesternight's 1 unlike 1 danger. 1 lips, 1 pretence 1 seized. 1 deferred 1 visit. 1 replaced 1 teachers 1 Besides, 1 nonsense?" 1 life. 1 guide 1 promised 1 secluded 1 inquirers 1 almost 1 engaged 1 study; 1 destiny. 1 You 1 arrive, 1 seem 1 watchful 1 away, 1 erroneously 1 fate 1 seeking 1 imbued 1 "I 1 who 1 you," 1 arguments 1 deference 1 stepped 1 disciple 1 grandeur 1 Alas! 1 arrives 1 scarcely 1 commenced, 1 evil 1 moment 1 transmuted 1 student 1 been, 1 palpable 1 events, 1 laboratory 1 totally 1 greedily 1 enchanting 1 event. 1 studied. 1 shortly 1 chimera 1 asked 1 person 1 expected, 1 exhibited. 1 unfitted 1 spend 1 left 1 benignity 1 idleness 1 endeavour 1 departed 1 less 1 indulge 1 removed 1 fancying 1 rest 1 ideas 1 schools 1 professor's 1 instructor, 1 affirmative. 1 facts 1 retired 1 happiness 1 myself. 1 letting 1 grappling 1 temples, 1 death 1 enthusiasm 1 experimentalist, 1 conclusions 1 alternate 1 shape. 1 pronouncing 1 parents 1 attractive 1 derange 1 Destruction, 1 By 1 minute," 1 read 1 room, 1 unlimited 1 know 1 destroy 1 press 1 dreams 1 preparatory 1 dignity 1 earthquake, 1 necessary 1 contempt, 1 after. 1 marked, 1 enounced 1 country. 1 zeal. 1 zeal 1 continue 1 chemist 1 view 1 works 1 inclined 1 worth. 1 vain. 1 old 1 often 1 requested 1 "promised 1 back 1 dream. 1 fifty 1 sight 1 done, 1 home 1 menaced, 1 "The 1 apply 1 pioneer 1 cooped 1 content 1 commences. 1 scientific 1 power 1 Geneva, 1 procure 1 disappointed, 1 respite 1 father. 1 preserver. 1 Chemistry 1 forget. 1 about 1 actual 1 visions 1 pleased. 1 hiding-places. 1 urged 1 despair 1 carelessly, 1 severe, 1 memorable 1 countenance; 1 desires 1 chimeras 1 letters 1 smiled 1 Magnus 1 instruments 1 talent. 1 down 1 education. 1 promise 1 narration 1 names. 1 endeavours 1 dirt, 1 endeavouring 1 assumed 1 restrained 1 Paracelsus, 1 Paracelsus. 1 much 1 happy 1 head 1 insurrection 1 form 1 imbibed 1 becoming 1 dabble 1 philosophers 1 malignity 1 anew." 1 you; 1 prognosticated 1 children. 1 being; 1 ear 1 deepest 1 also 1 rush 1 veiled 1 chained 1 invincible 1 mechanism. 1 necessity; 1 up 1 placed 1 carriage 1 limit 1 home, 1 he, 1 eyes. 1 alarm 1 affection 1 advise 1 friend. 1 liberal 1 pore 1 certain 1 Ingolstadt. 1 lost. 1 metals 1 scarlet 1 proves 1 ensuing 1 student, 1 education 1 internal 1 mutual 1 mankind." 1 philosophy, 1 Never 1 mimic 1 reality 1 application 1 details 1 department 1 unwilling 1 residence 1 lectures. 1 mock 1 smiles 1 ancient? 1 formed 1 impossibilities 1 "Have 1 indeed, 1 favourite 1 omen, 1 ultimately 1 resign 1 town 1 deathbed 1 sir, 1 utterly 1 death, 1 death. 1 friends 1 died 1 omnipotent 1 turmoil; 1 younger 1 land 1 longer 1 recapitulation 1 age 1 required 1 rose. 1 conception, 1 longed 1 At 1 treading 1 resolution 1 having 1 once 1 