the 134 of 114 and 95 to 75 my 51 I 50 a 46 was 41 in 33 that 24 with 24 were 19 which 17 by 15 had 15 but 14 not 12 for 12 from 11 our 11 their 11 as 11 this 10 it 10 we 9 It 9 me 8 so 8 have 8 he 8 all 7 spirit 7 its 7 his 7 He 7 on 7 or 7 an 7 When 6 The 6 her 6 at 6 even 5 My 5 more 5 they 5 could 5 are 5 those 5 myself 5 upon 5 into 5 father 4 would 4 soul 4 than 4 most 4 We 4 been 4 is 4 studies. 4 if 4 possessed 4 like 4 up 4 seemed 3 science 3 me. 3 nature, 3 while 3 new 3 men 3 great 3 changed 3 former 3 man 3 always 3 entirely 3 house 3 philosophy 3 one 3 such 3 was, 3 natural 3 occupied 3 laws 3 soon 3 she 3 secrets 3 Cornelius 3 among 3 life 3 mind 3 these 3 might 3 never 3 greatest 3 In 3 human 3 but, 3 parents 3 real 3 read 3 acquainted 3 beheld 3 Clerval 3 own 3 there 3 us 3 knowledge. 3 once 3 very 2 more. 2 me, 2 deeply 2 ever 2 led 2 ruin. 2 desired 2 myself. 2 glance 2 should 2 thus 2 train 2 effort 2 learn 2 Belrive, 2 discovery 2 terrible 2 rather 2 stood 2 singular 2 All 2 light 2 tale 2 pleasure 2 years 2 still 2 powers 2 greater 2 She 2 kindness 2 adventurous 2 nor 2 found 2 therefore, 2 Elizabeth 2 thirst 2 research 2 theory 2 wonderful 2 passed 2 exploded 2 modern 2 Albertus 2 any 2 latter 2 subject 2 who 2 storm 2 find 2 about 2 various 2 him 2 violent 2 gladness 2 said 2 here 2 many 2 became 2 afterwards 2 Her 2 appeared 2 unfolded 2 entered 2 And 2 delight. 2 near 2 Agrippa 2 almost 2 engaged 2 things 2 ardour 2 characters 2 being 2 oak 2 facts 2 followed 2 taken 2 has 2 gave 2 On 2 early 2 birth 2 become 2 works 2 old 2 home 2 passion 2 be 2 knew 2 Geneva, 2 intense 2 utterly 2 nothing 2 But 2 lot 2 some 2 volume 2 made 2 temper 2 when 2 favourite 2 felt 2 time 2 childish 2  1 code 1 impulse 1 son, 1 branches 1 soften 1 thoughtful 1 philosopher 1 hanging 1 ignorantly 1 causes 1 whose 1 certainly 1 fancies 1 catastrophe, 1 seems 1 tranquillity 1 under 1 carelessly 1 immutable 1 Nor 1 merchant 1 cause, 1 attempts 1 returned 1 returning 1 rashly 1 wood. 1 souls 1 gloomy 1 Henry 1 theme; 1 word 1 difference 1 continued 1 busied 1 heaven 1 went 1 sought; 1 knightly 1 tenderness 1 progress 1 disciple. 1 frightful 1 inclination 1 added 1 deformed 1 object, 1 decreed 1 indifferent, 1 second 1 entertained 1 utter 1 ardent 1 desire, 1 tempest 1 penetrated 1 lineaments 1 what 1 plays 1 appear 1 Agrippa. 1 witnessed 1 assisted 1 general; 1 Clerval? 1 him. 1 century; 1 then 1 unadept, 1 learned 1 contrast 1 thin 1 full 1 avert 1 guardian 1 languages, 1 drew 1 river, 1 will 1 yards 1 imagination; 1 strong 1 change 1 obtained 1 boy 1 substance 1 talent 1 study 1 electricity 1 within 1 principally 1 narrow 1 changes 1 guidance 1 composed 1 love 1 danger 1 suddenly 1 retired 1 elixir 1 brought 1 vanished, 1 moral 1 names 1 Isaac 1 tertiary 1 untaught 1 give 1 beneficence 1 few 1 circumstances 1 warmed 1 mysterious 1 scope 1 themselves 1 liberally 1 burst 1 Those 1 holy 1 instructors. 1 apprehensions 1 known 1 companionship, 1 violent, 1 mountains 1 shrine-dedicated 1 account 1 fatal 1 avidity. 1 us. 1 us, 1 imagination, 1 theories 1 himself, 1 remain 1 sudden 1 obvious 1 can 1 following 1 akin 1 history 1 beautiful 1 lords 1 want 1 stream 1 baths 1 shattered 1 states 1 inexperience 1 unveiled 1 arise 1 cursory 1 species 1 galvanism, 1 native 1 summers 1 attract; 1 united 1 end 1 ideas 1 means 1 fortunate 1 write 1 how 1 lamp 1 writers 1 youth, 1 degree, 1 steps, 1 entrench 1 A 1 systems, 1 tried 1 attend 1 may 1 fancy. 1 after 1 stars 1 blood 1 blindness, 1 accorded 1 Swiss 1 waste 1 heroes 1 law 1 tormenting 1 abortive 1 introduced 1 speak, 1 averred, 1 fortifications 1 shore 1 shade 1 enter 1 calm, 1 dream 1 make 1 Thonon; 1 satisfied 1 bounding 1 known. 1 through 1 gazed 1 fidelity 1 inquiries 1 before 1 till 1 progeny 1 inferior 1 course, 1 gentleness. 1 author, 1 creations 1 whole 1 subsisted 1 hidden 1 world. 1 led, 1 pursue 1 good 1 tyrants 1 ancient, 1 ineffectual. 1 names; 1 thirteen 1 recollections 1 hands 1 desperately 1 constructed, 1 Newton 1 creation, 1 bless 1 peasant 1 victory 1 each 1 predilection 1 friendship 1 potent, 1 exquisite 1 Magnus, 1 bright 1 Destiny 1 doing 1 pursuits 1 dispute. 1 books 1 Harmony 1 entering 1 year 1 dawn 1 gallant 1 living 1 misfortune 1 mind, 1 confess 1 surrounded 1 despicable. 1 strangers 1 wondrous 1 current 1 issue 1 announced 1 Alpine 1 appertaining 1 unacquainted 1 assured 1 associate 1 title 1 envelop 1 little 1 quite 1 pursuit. 1 struggle 1 besides 1 earliest 1 heroic 1 care 1 thrown 1 attention. 1 things. 1 relinquishing 1 things, 1 overthrow 1 contented 1 keep 1 inclemency 1 sensations 1 twenty 1 loudness 1 childhood 1 first 1 Victor, 1 chimerical, 1 Agrippa, 1 dwelling 1 curiosity 1 render 1 Jura, 1 feel 1 attractions 1 preservation 1 sympathy 1 soaring 1 Roncesvalles, 1 long 1 generosity, 1 If, 1 filial 1 visions 1 remember. 1 story 1 ancient 1 temperature 1 attach 1 families 1 unknown 1 love. 1 system 1 relations 1 too 1 perfectly 1 final 1 boy's 1 disposition; 1 pains 1 explanation 1 studies 1 took 1 immediate 1 treasures 1 repined. 1 herself 1 loved 1 grew 1 aught 1 joys. 1 scenes 1 heavens. 1 visited 1 seclusion. 1 wandering 1 torrent 1 sublime 1 usefulness 1 metaphysical, 1 hardship, 1 angel 1 remark, 1 chivalrous 1 disunion 1 turned 1 sad 1 threw 1 say 1 need 1 saintly 1 secure 1 built 1 diligence 1 aside 1 eagerly 1 preceptors 1 also 1 labour 1 invulnerable 1 towards 1 student's 1 procure 1 voice, 1 disappeared, 1 thunder 1 childhood, 1 bound 1 indiscriminately. 1 failure 1 door, 1 sometimes 1 science. 1 disease 1 face 1 looked 1 sepulchre 1 "Ah! 1 reflections 1 Agrippa! 1 tainted 1 nature. 1 came 1 occupations, 1 regulated 1 swelling 1 proceeded, 1 indulgence. 1 ardour, 1 Under 1 threshold 1 earth 1 rough 1 chanced 1 nearer 1 busy 1 spite 1 Meanwhile 1 poets; 1 consideration. 1 explain 1 behind 1 worthy 1 considerable 1 unsuccessful, 1 incantations 1 only 1 watching 1 partially 1 few. 1 guided 1 hope 1 do 1 bonds 1 remained, 1 While 1 vehement; 1 foundations, 1 distinctly 1 penetrate 1 quarters 1 tyros 1 secondary 1 glory 1 contents, 1 species. 1 them. 1 fixed 1 communicated 1 insensible 1 caprice, 1 loveliness 1 set 1 city. 1 Wealth 1 swept 1 devils 1 tree 1 frame 1 eighteenth 1 Paracelsus 1 trash." 1 outward 1 wonder 1 destiny 1 caprices 1 study, 1 self-taught 1 away 1 adventure. 1 genius 1 state 1 ages. 1 years, 1 routine 1 drawn 1 neither 1 heroes, 1 King 1 romance. 1 Natural 1 nature 1 attention 1 ideas. 1 days, 1 infidels. 1 floundering 1 fatality 1 inn. 1 picking 1 blasted 1 concentrated 1 league 1 feeling 1 last 1 disdain 1 ill 1 learn; 1 according 1 attributed 1 resided 1 prosecution, 1 joy, 1 forgotten 1 ambition. 1 learn, 1 Yet 1 masquerades, 1 together; 1 impediments 1 Sir 1 sweet 1 winter, 1 enterprise, 1 Nature, 1 agents 1 together. 1 majestic 1 reasoning, 1 sense, 1 speak 1 gratitude 1 unusual 1 described 1 capable 1 fifteen 1 remained 1 dazzling 1 whom 1 secret 1 much 1 philosophers, 1 peaceful 1 apathy; 1 home. 1 delights 1 citadel 1 shock, 1 diversity 1 deeper 1 eastern 1 fire 1 thousand 1 formed 1 search 1 manner. 1 accident 1 lives 1 child 1 uses. 1 Round 1 banish 1 look 1 contemplated 1 life; 1 By 1 aim 1 delight; 1 Besides, 1 wild 1 investigating 1 life, 1 discoveries 1 mistake 1 seven 1 studied 1 ligaments 1 lasted, 1 unsatisfied. 1 ready 1 said, 1 dissect, 1 would-be 1 perhaps 1 began 1 imbued 1 same 1 beside 1 strange 1 disregard. 1 party 1 immortal 1 events 1 day 1 development 1 noble 1 suggestion 1 closest 1 mountain 1 rapture, 1 appearances 1 evil 1 companion 1 authors, 1 Curiosity, 1 governments, 1 longing 1 successors 1 narration, 1 no 1 ocean 1 which, 1 Table 1 creators 1 drawing 1 betook 1 left 1 scientific, 1 actions 1 ignoble 1 schools 1 grades 1 turbulence 1 skill 1 happiness 1 undivided 1 latter, 1 eager 1 book 1 destruction. 1 visions. 1 extensive 1 excited 1 around 1 ample 1 possible 1 practical, 1 earnest 1 redeem 1 truth. 1 confined 1 world 1 exploit, 1 advanced 1 ruled 1 desire 1 causes. 1 country. 1 multifarious 1 shapes 1 miraculous 1 campagne 1 soft 1 page 1 Before 1 unexplored 1 shed 1 because 1 crowd 1 obliged 1 magnificent 1 disinclined 1 humane, 1 lake, 1 elements 1 dear 1 animate 1 passions 1 mood 1 arise, 1 avoid 1 recorded 1 shone 1 sake. 1 good, 1 slight 1 Geneva. 1 peculiarly 1 virtues 1 destroyed. 1 step 1 mystery. 1 calmer 1 father. 1 stage 1 stone 1 discontented 1 mingled 1 anything 1 enjoyed. 1 reduced 1 practical 1 greatly 1 act 1 self. 1 benefactors 1 silence 1 chivalry 1 No 1 electricity. 1 delighted 1 son 1 down 1 beings 1 weather 1 promise 1 mingling, 1 next 1 morning, 1 your 1 anatomize, 1 strangely 1 shells 1 splintered 1 amidst 1 fervent 1 Paracelsus, 1 avowed 1 inner 1 seasons, 1 prosperity 1 books, 1 slough 1 child's 1 enchantment 1 regard 1 principles 1 misery, 1 contradictory 1 Arthur, 1 hopes 1 highest 1 junior 1 raising 1 directed 1 admiration 1 philosopher's 1 whether 1 Magnus. 1 record 1 taught 1 accustomed 1 divine. 1 fate; 1 demonstrate 1 this; 1 eyes, 1 enthusiasm. 1 distance 1 instead 1 celestial 1 aerial 1 subdue 1 house; 1 received 1 imagination 1 relates 1 politics 1 education 1 ghosts 1 smile, 1 physical 1 again 1 knowledge, 1 sullen 1 sources; 1 astonishing 1 discerned 1 back, 1 application 1 other 1 branch 1 latterly 1 mathematics 1 thunderstorm. 1 ribbons 1 picture 1 semblance 1 smitten 1 ours; 1 death! 1 fervently 1 occasion 1 structure 1 opened 1 school-fellows 1 happier 1 age 1 stump. 1 Thus 1 rule 1 having 1 As 1 serious 1 fulfilment 1 mountains, 1 songs 1 