of 74 and 69 the 68 to 61 a 52 her 42 was 39 in 32 my 29 his 27 had 24 their 20 that 16 by 15 he 15 with 13 for 12 on 12 father 11 it 11 I 11 she 10 as 10 but 10 from 9 they 9 all 8 this 8 which 8 one 7 The 7 He 7 seemed 6 years 6 than 6 became 6 Her 6 mother 6 been 6 while 5 more 5 so 5 him 5 them 5 She 5 were 5 an 5 when 5 me 4 My 4 not 4 could 4 mine 4 who 4 only 4 Beaufort 4 child 4 being 4 be 4 at 4 whose 3 mother, 3 very 3 child, 3 benevolent 3 me. 3 what 3 public 3 poverty 3 daughter 3 after 3 infant 3 through 3 There 3 little 3 passed 3 mind 3 have 3 most 3 means 3 these 3 They 3 some 3 months 3 made 3 no 3 died 3 Elizabeth 3 time 3 attracted 2 pride 2 eldest 2 every 2 Milan, 2 her. 2 her, 2 During 2 love 2 When 2 charge 2 found 2 circumstances 2 attachment 2 creature 2 One 2 His 2 continued 2 name 2 peasant 2 each 2 accompanied 2 Caroline 2 beggar. 2 This 2 disposition 2 Italy, 2 long 2 friend 2 eyes 2 loved 2 marriage 2 visited 2 distinguished 2 With 2 towards 2 its 2 I, 2 abode. 2 during 2 yield 2 them. 2 where 2 set 2 orphan 2 father's 2 girl, 2 received 2 rose 2 But 2 life 2 sufficient 2 spirit 2 Italy 2 is 2 fairer 2 occupied 2 several 2 upon 2 among 2 previous 2 five 2 about 2 despair 2 or 2 support 2 there 2 himself 2 placed 2 affection 2 gone 2 deep 2 other 2 better 2 poor 2 bestowed 2  1 Reuss. 1 knelt 1 month 1 four 1 integrity 1 children 1 devoted 1 praises 1 former 1 duty; 1 foster 1 those 1 tranquillity 1 under 1 smile 1 suffered 1 merchant 1 garden 1 wretchedness. 1 wishes 1 emotion 1 difference 1 child. 1 poor. 1 singularly 1 tenderness 1 small 1 moulding 1 added 1 ten 1 other, 1 me, 1 direct 1 street 1 honourable 1 helpless 1 expressive 1 situated 1 even 1 pittance 1 mould, 1 wreck 1 giving 1 saved 1 sum 1 liberty 1 gold, 1 him. 1 prevailed 1 rest. 1 above 1 conduct 1 filled 1 strongly. 1 body 1 led 1 honour 1 gathered 1 vale 1 behaviour 1 desired 1 entered, 1 same 1 alone 1 change 1 through. 1 animated 1 bloomed 1 inspired 1 leaving 1 credit 1 cherish. 1 misery 1 sweetness 1 worse; 1 Victor 1 family 1 straw 1 inexhaustible 1 highly 1 sorrows 1 hardy 1 chamois 1 spoke 1 would 1 sister, 1 two 1 distributing 1 live 1 suffered, 1 shaken 1 weeping 1 bitterly 1 taken 1 until 1 possession 1 pretty 1 evening 1 subsistence 1 orphan. 1 wonders, 1 sister 1 refrain 1 grief 1 train 1 bitterly, 1 hold 1 town 1 none 1 hour 1 retreated 1 himself, 1 thin 1 making 1 coffin 1 lingered 1 beautiful 1 German 1 radiance 1 self-control, 1 bent 1 gardener, 1 convenience. 1 offspring. 1 endured, 1 something 1 want 1 sense 1 sought 1 clothing, 1 Several 1 deplored 1 returned 1 united 1 end 1 provide 1 bonds 1 conducted 1 how 1 procured 1 Beaufort's 1 frontiers 1 confiscated; 1 relinquished 1 Their 1 playfully, 1 assistance. 1 protection 1 may 1 state, 1 shores 1 ample, 1 bear 1 vagrants; 1 contrived 1 All 1 Everyone 1 consulted 1 France. 1 courage 1 decreasing 1 wife, 1 pleasure 1 first 1 words 1 playing 1 wind 1 affection. 1 lighter 1 idol, 1 welcomed 1 unworthiness 1 soon 1 strove 1 early, 1 motions 1 committed 1 still 1 worship 1 before 1 rapidly 1 Overjoyed 1 till 1 No 1 months, 1 fair. 1 meantime 1 pleasurable 1 married, 1 truest 1 greater 1 indefatigable 1 regarding 1 history. 1 number 1 hands 1 hitherto 1 hall 1 nor 1 frementi, 1 Everything 1 degree, 1 labour, 1 entirely 1 friendship 1 meal 1 mean 1 afforded 1 From 1 scanty 1 house 1 hard 1 house. 1 house, 1 health, 1 therefore, 1 our 1 tenth 1 event 1 brow 1 tried 1 decreased; 1 overcame 1 both, 1 childish 1 since 1 wholly 1 looking 1 enjoyment 1 day, 1 features. 1 forth 1 attended 1 circumstance 1 given 1 pleasant 1 attending 1 bestow 1 born. 1 brightest 1 attendant 1 care 1 support. 1 them, 1 persuading 1 days 1 protection. 1 keep 1 turn 1 length 1 familiarly 1 family. 1 lay 1 exotic 1 syndics, 1 occupations 1 sickness, 1 dungeons 1 powerful 1 scene 1 rank 1 such 1 tomorrow 1 illustrate 1 Elizabeth. 1 abode, 1 For 1 unknown 1 inmate 1 relieved 1 morrow, 1 took 1 inexpressible 1 was, 1 of, 1 love, 1 herself 1 grace 1 disconsolate, 1 reverential 1 grew 1 fell, 1 bed 1 relation. 1 exertion. 1 prospect 1 false 1 angel 1 remained 1 saw 1 any 1 affairs 1 cottages 1 reflection, 1 patience, 1 Germany 1 blue 1 begin 1 beyond 1 shall 1 procure 1 paid 1 This, 1 age, 1 reverence 1 inaction; 1 stood 1 future 1 him; 1 afflicted. 1 clear 1 proud 1 hungry 1 face 1 looked 1 perceiving 1 deeply 1 came 1 penury 1 show 1 word, 1 fond 1 reputation. 1 discovered 1 bring 1 relation 1 imagined 1 debts, 1 We 1 just 1 justice 1 situations 1 should 1 mind. 1 plaited 1 excursion 1 priest, 1 hope 1 heaven, 1 Whether 1 kind 1 leisure 1 unfair 1 cannot 1 circumstances. 1 despite 1 interpreted 1 Having 1 stamp 1 earn 1 late-discovered 1 numerous 1 doting 1 seriousness, 1 effectual 1 cousin. 1 fixed 1 communicated 1 husband 1 looks 1 victim 1 fair 1 exerted 1 are 1 rankling 1 tender 1 hastened 1 wonder 1 closer 1 said 1 tend 1 various 1 between 1 promised 1 man, 1 notice 1 chamber. 1 dark-leaved 1 attention 1 antique 1 Genevese, 1 unbending 1 rude 1 head. 1 then. 1 grieved 1 climate 1 necessity, 1 last 1 cot 1 when, 1 rambles. 1 many 1 according 1 old, 1 fulfilled 1 adored 1 tour 1 present 1 distinction 1 spirit, 1 approve 1 pleasures. 1 bearing 1 appeared 1 charity, 1 others 1 active 1 foldings 1 village 1 constant 1 rougher 1 poverty. 1 gratitude 1 decline 1 union 1 own. 1 three 1 whom 1 much 1 interest 1 became, 1 entered 1 lovely 1 duties 1 lived 1 innocent 1 Among 1 ages 1 blessing 1 excite 1 uncommon 1 manner. 1 fund 1 manner, 1 protect, 1 mischances, 1 Lucerne, 1 And 1 delight. 1 plain 1 value 1 care; 1 who, 1 near 1 parents' 1 country 1 life. 1 care. 1 life, 1 parents, 1 known. 1 remembering 1 owed 1 working, 1 almost 1 character, 1 sustenance 1 respected 1 birth. 1 good 1 property 1 result 1 different 1 consequently, 1 perpetually 1 "I 1 unite 1 it." 1 prevented 1 sheltered 1 unfortunate 1 heaven-sent, 1 week 1 differing 1 companion 1 guardians 1 guardian 1 cherub 1 single 1 nobleman. 1 villa 1 daughter, 1 scarcely 1 off 1 weakened 1 mother's 1 expression 1 possessed 1 variety 1 spent 1 dark-eyed, 1 babes. 1 without 1 greatest 1 incapable 1 schiavi 1 stores 1 consciousness 1 money 1 guided 1 obtain 1 republic. 1 eagerly 1 tenderness, 1 immediately 1 protecting 1 happiness 1 blow 1 death 1 apparition 1 marrying 1 regarded 1 brambles. 1 shape. 1 knew 1 work; 1 parents 1 beloved 1 sweet 1 gift, 1 Como. 1 gave 1 silken 1 On 1 wife. 1 elapsed 1 birth 1 world 1 behold 1 retreat 1 desire 1 brought 1 necessary 1 like 1 lost 1 Providence 1 seek 1 country. 1 cloudless, 1 oblivion 1 counsellors 1 country; 1 passionate 1 soft 1 half-clothed 1 worth. 1 shed 1 often 1 people 1 it, 1 hair 1 born 1 lips 1 Much 1 interment 1 employment 1 gradually 1 literally 1 passion 1 flourishing 1 good, 1 cord 1 measures 1 merchant's 1 intimate 1 virtues 1 business. 1 woman, 1 worthy 1 weakness. 1 relating 1 fondness 1 conceal 1 ognor 1 surround 1 distinct 1 Austria 1 act 1 shared 1 permission 1 out, 1 enter 1 adversity. 1 rendered 1 restorative 1 formerly 1 presence 1 into 1 Two 1 down 1 respectable 1 lesson 1 rustic 1 endeavouring 1 disposed 1 fast 1 only. 1 caresses 1 lot 1 worst 1 recollections. 1 hills. 1 Lavenza 1 frame. 1 form 1 crown 1 memory 1 hoped 1 misery, 1 upright 1 Italians 1 considerable 1 admiration 1 glory 1 species, 1 fortunes, 1 attached 1 up 1 home, 1 plaything 1 called 1 celestial 1 discovery, 1 stock. 1 Beaufort, 1 Perhaps 1 am 1 Lake 1 arms, 1 walks 1 nursed 1 again 1 explained. 1 ancestors 1 Geneva 1 magnificence. 1 Milanese 1 Naples, 1 nurse: 1 draw 1 living 1 shelter 1 recompensing 1 friends 1 younger 1 land 1 interval 1 pictured 1 functions; 1 As 1 presented 1 far 1 sensibility 1 